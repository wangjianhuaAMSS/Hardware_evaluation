module M(f_in, f_out);
    input [63 : 0] f_in;
    output [63: 0] f_out;
      assign f_out[63] = f_in[59] ^ f_in[55] ^ f_in[51];
      assign f_out[62] = f_in[62] ^ f_in[54] ^ f_in[50];
      assign f_out[61] = f_in[61] ^ f_in[57] ^ f_in[49];
      assign f_out[60] = f_in[60] ^ f_in[56] ^ f_in[52];
      assign f_out[59] = f_in[63] ^ f_in[59] ^ f_in[55];
      assign f_out[58] = f_in[58] ^ f_in[54] ^ f_in[50];
      assign f_out[57] = f_in[61] ^ f_in[53] ^ f_in[49];
      assign f_out[56] = f_in[60] ^ f_in[56] ^ f_in[48];
      assign f_out[55] = f_in[63] ^ f_in[59] ^ f_in[51];
      assign f_out[54] = f_in[62] ^ f_in[58] ^ f_in[54];
      assign f_out[53] = f_in[57] ^ f_in[53] ^ f_in[49];
      assign f_out[52] = f_in[60] ^ f_in[52] ^ f_in[48];
      assign f_out[51] = f_in[63] ^ f_in[55] ^ f_in[51];
      assign f_out[50] = f_in[62] ^ f_in[58] ^ f_in[50];
      assign f_out[49] = f_in[61] ^ f_in[57] ^ f_in[53];
      assign f_out[48] = f_in[56] ^ f_in[52] ^ f_in[48];
      assign f_out[47] = f_in[47] ^ f_in[43] ^ f_in[39];
      assign f_out[46] = f_in[42] ^ f_in[38] ^ f_in[34];
      assign f_out[45] = f_in[45] ^ f_in[37] ^ f_in[33];
      assign f_out[44] = f_in[44] ^ f_in[40] ^ f_in[32];
      assign f_out[43] = f_in[47] ^ f_in[43] ^ f_in[35];
      assign f_out[42] = f_in[46] ^ f_in[42] ^ f_in[38];
      assign f_out[41] = f_in[41] ^ f_in[37] ^ f_in[33];
      assign f_out[40] = f_in[44] ^ f_in[36] ^ f_in[32];
      assign f_out[39] = f_in[47] ^ f_in[39] ^ f_in[35];
      assign f_out[38] = f_in[46] ^ f_in[42] ^ f_in[34];
      assign f_out[37] = f_in[45] ^ f_in[41] ^ f_in[37];
      assign f_out[36] = f_in[40] ^ f_in[36] ^ f_in[32];
      assign f_out[35] = f_in[43] ^ f_in[39] ^ f_in[35];
      assign f_out[34] = f_in[46] ^ f_in[38] ^ f_in[34];
      assign f_out[33] = f_in[45] ^ f_in[41] ^ f_in[33];
      assign f_out[32] = f_in[44] ^ f_in[40] ^ f_in[36];
      assign f_out[31] = f_in[31] ^ f_in[27] ^ f_in[23];
      assign f_out[30] = f_in[26] ^ f_in[22] ^ f_in[18];
      assign f_out[29] = f_in[29] ^ f_in[21] ^ f_in[17];
      assign f_out[28] = f_in[28] ^ f_in[24] ^ f_in[16];
      assign f_out[27] = f_in[31] ^ f_in[27] ^ f_in[19];
      assign f_out[26] = f_in[30] ^ f_in[26] ^ f_in[22];
      assign f_out[25] = f_in[25] ^ f_in[21] ^ f_in[17];
      assign f_out[24] = f_in[28] ^ f_in[20] ^ f_in[16];
      assign f_out[23] = f_in[31] ^ f_in[23] ^ f_in[19];
      assign f_out[22] = f_in[30] ^ f_in[26] ^ f_in[18];
      assign f_out[21] = f_in[29] ^ f_in[25] ^ f_in[21];
      assign f_out[20] = f_in[24] ^ f_in[20] ^ f_in[16];
      assign f_out[19] = f_in[27] ^ f_in[23] ^ f_in[19];
      assign f_out[18] = f_in[30] ^ f_in[22] ^ f_in[18];
      assign f_out[17] = f_in[29] ^ f_in[25] ^ f_in[17];
      assign f_out[16] = f_in[28] ^ f_in[24] ^ f_in[20];
      assign f_out[15] = f_in[11] ^ f_in[07] ^ f_in[03];
      assign f_out[14] = f_in[14] ^ f_in[06] ^ f_in[02];
      assign f_out[13] = f_in[13] ^ f_in[09] ^ f_in[01];
      assign f_out[12] = f_in[12] ^ f_in[08] ^ f_in[04];
      assign f_out[11] = f_in[15] ^ f_in[11] ^ f_in[07];
      assign f_out[10] = f_in[10] ^ f_in[06] ^ f_in[02];
      assign f_out[09] = f_in[13] ^ f_in[05] ^ f_in[01];
      assign f_out[08] = f_in[12] ^ f_in[08] ^ f_in[00];
      assign f_out[07] = f_in[15] ^ f_in[11] ^ f_in[03];
      assign f_out[06] = f_in[14] ^ f_in[10] ^ f_in[06];
      assign f_out[05] = f_in[09] ^ f_in[05] ^ f_in[01];
      assign f_out[04] = f_in[12] ^ f_in[04] ^ f_in[00];
      assign f_out[03] = f_in[15] ^ f_in[07] ^ f_in[03];
      assign f_out[02] = f_in[14] ^ f_in[10] ^ f_in[02];
      assign f_out[01] = f_in[13] ^ f_in[09] ^ f_in[05];
      assign f_out[00] = f_in[08] ^ f_in[04] ^ f_in[00];

endmodule